module MUX2_1();
endmodule
